`include "opcodes.v"

module CPU (
  output [31:0] pc,
  input         clk,
  input  [31:0] instruction
);
endmodule
