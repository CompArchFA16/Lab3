`ifndef __MUX_T_V__
`define __MUX_T_V__
module test_mux();

initial begin

end

endmodule
`endif
