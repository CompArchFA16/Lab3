// TODO: Move these tests into the main file after we consolidate.

module testDavidsStuff ();

  initial begin

    // J =======================================================================

    // JR ======================================================================

    // JAL =====================================================================

    // JSUB ====================================================================

  end
endmodule
