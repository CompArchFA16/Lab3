`include "opcodes.v"
`include "gate_ID_EX.v"

module CPU (
  output [31:0] pc,
  input         clk,
  input  [31:0] instruction
);
endmodule
